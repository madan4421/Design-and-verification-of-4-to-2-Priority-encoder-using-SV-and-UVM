interface pe_interface();
    logic [3:0] in;
    logic [1:0] out;
    logic valid;     
endinterface  